module and2(Y, A, B);
	input A, B;
	output Y;
	and (Y, A, B);
endmodule