library verilog;
use verilog.vl_types.all;
entity and2_tb is
end and2_tb;
